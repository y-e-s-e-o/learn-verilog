module not_gate(A_i, F_o);
    
    input A_i;
    output F_o;
    assign F_o = ~A_i;

endmodule